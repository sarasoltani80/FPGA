
module correlation_32_tb;

reg [31:0] Num_1, Num_2, Num_3, Num_4, Num_5, Num_6, Num_7, Num_8, Num_9, Num_10, Num_11, Num_12, Num_13, Num_14, Num_15, Num_16,  Target_Num;
reg Clock, Reset;

wire [3:0] out_4;

  correlation_32 u (Num_1, Num_2, Num_3, Num_4, Num_5, Num_6, Num_7, Num_8, Num_9, Num_10, Num_11, Num_12, Num_13, Num_14, Num_15, Num_16,Target_Num,Clock,Reset,out_4);

  initial begin

    Clock = 0;
    Reset = 1;
    Num_1 = 32'b0;
    Num_2 = 32'b0;
    Num_3 = 32'b0;
    Num_4 = 32'b0;
    Num_5 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_6 = 32'b0;
    Num_7 = 32'b0;
    Num_8 = 32'b0;
    Num_9 = 32'b0;
    Num_10 = 32'b0;
    Num_11 = 32'b0;
    Num_12 = 32'b0;
    Num_13 = 32'b0;
    Num_14 = 32'b0;
    Num_15 = 32'b0;
    Num_16 = 32'b0;
    Target_Num = 32'b1111_1111_1111_1111_1111_1111_1111_1111;

$monitor("%d  Clock=%b, Reset=%b, Num_1=%b, Num_2=%b, Num_3=%b, Num_4=%b, Num_5=%b, Num_6=%b, Num_7=%b, Num_8=%b, Num_9=%b, Num_10=%b, Num_11=%b, Num_12=%b, Num_13=%b, Num_14=%b, Num_15=%b, Num_16=%b, Target_Num=%b, out_4=%b",$time,
 Clock, Reset, Num_1, Num_2, Num_3, Num_4, Num_5, Num_6, Num_7, Num_8, Num_9, Num_10, Num_11, Num_12, Num_13, Num_14, Num_15, Num_16,  Target_Num, out_4);


  #5;
     Num_1 = 32'b0;
    Num_2 = 32'b0;
    Num_3 = 32'b0;
    Num_4 = 32'b0;
    Num_5 = 32'b0;
    Num_6 = 32'b0;
    Num_7 = 32'b0;
    Num_8 = 32'b0;
    Num_9 = 32'b0;
    Num_10 = 32'b0;
    Num_11 = 32'b0;
    Num_12 = 32'b0;
    Num_13 = 32'b0;
    Num_14 = 32'b0;
    Num_15 = 32'b0;
    Num_16 = 32'b0;
    Reset=0;

    #10;
    Num_1 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_3 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_4 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_16 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
#5 Reset=1;

    #10;
Reset=0;
    Num_2 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_3 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_4 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_16 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

   #10;
    Num_3 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_4 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_16 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

    #10;
    Num_4 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_3 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_16 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

   #10;
    Num_4 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_3 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b1111_1111_1111_1111_1111_1111_1111_1100;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b1111_1111_1111_1000_1111_1111_1111_1111;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_16 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

   #10;
    Num_16 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_3 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_4 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

   #10;
    Num_4 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Num_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_3 = 32'b1111_1001_1111_1111_1111_1111_1111_1100; 
    Num_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_5 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_6 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_7 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_8 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_9 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_10 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_11 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_12 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_13 = 332'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_14 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_15 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Num_16 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

    
  end
  initial repeat (20) #5 Clock = ~Clock;

endmodule

